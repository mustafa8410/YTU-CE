module zeroExtend_1bit(a,out);
    input a;
    output out;
    assign out = a;
endmodule